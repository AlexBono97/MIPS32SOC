//  A testbench for testMemoryRDataDecoder_tb
`timescale 1us/1ns

module testMemoryRDataDecoder_tb;
    reg [31:0] dIn;
    reg [1:0] offset;
    reg dExt;
    reg [1:0] dSize;
    wire [31:0] dOut;

  testMemoryRDataDecoder testMemoryRDataDecoder0 (
    .dIn(dIn),
    .offset(offset),
    .dExt(dExt),
    .dSize(dSize),
    .dOut(dOut)
  );

    reg [68:0] patterns[0:23];
    integer i;

    initial begin
      patterns[0] = 69'b10101010101110111100110011011101_00_0_00_10101010101110111100110011011101;
      patterns[1] = 69'b10101010101110111100110011011101_01_0_00_10101010101110111100110011011101;
      patterns[2] = 69'b10101010101110111100110011011101_10_0_00_10101010101110111100110011011101;
      patterns[3] = 69'b10101010101110111100110011011101_11_0_00_10101010101110111100110011011101;
      patterns[4] = 69'b10101010101110111100110011011101_00_1_00_10101010101110111100110011011101;
      patterns[5] = 69'b10101010101110111100110011011101_01_1_00_10101010101110111100110011011101;
      patterns[6] = 69'b10101010101110111100110011011101_10_1_00_10101010101110111100110011011101;
      patterns[7] = 69'b10101010101110111100110011011101_11_1_00_10101010101110111100110011011101;
      patterns[8] = 69'b10101010101110111100110011011101_00_0_01_00000000000000001010101010111011;
      patterns[9] = 69'b10101010101110111100110011011101_00_1_01_11111111111111111010101010111011;
      patterns[10] = 69'b10101010101110111100110011011101_01_0_01_00000000000000001010101010111011;
      patterns[11] = 69'b10101010101110111100110011011101_01_1_01_11111111111111111010101010111011;
      patterns[12] = 69'b10101010101110111100110011011101_10_0_01_00000000000000001100110011011101;
      patterns[13] = 69'b10101010101110111100110011011101_10_1_01_11111111111111111100110011011101;
      patterns[14] = 69'b10101010101110111100110011011101_11_0_01_00000000000000001100110011011101;
      patterns[15] = 69'b10101010101110111100110011011101_11_1_01_11111111111111111100110011011101;
      patterns[16] = 69'b10101010101110111100110011011101_00_0_10_00000000000000000000000010101010;
      patterns[17] = 69'b10101010101110111100110011011101_01_0_10_00000000000000000000000010111011;
      patterns[18] = 69'b10101010101110111100110011011101_10_0_10_00000000000000000000000011001100;
      patterns[19] = 69'b10101010101110111100110011011101_11_0_10_00000000000000000000000011011101;
      patterns[20] = 69'b10101010101110111100110011011101_00_1_10_11111111111111111111111110101010;
      patterns[21] = 69'b10101010101110111100110011011101_01_1_10_11111111111111111111111110111011;
      patterns[22] = 69'b10101010101110111100110011011101_10_1_10_11111111111111111111111111001100;
      patterns[23] = 69'b10101010101110111100110011011101_11_1_10_11111111111111111111111111011101;

      for (i = 0; i < 24; i = i + 1)
      begin
        dIn = patterns[i][68:37];
        offset = patterns[i][36:35];
        dExt = patterns[i][34];
        dSize = patterns[i][33:32];
        #10;
        if (patterns[i][31:0] !== 32'hx)
        begin
          if (dOut !== patterns[i][31:0])
          begin
            $display("%d:dOut: (assertion error). Expected %h, found %h", i, patterns[i][31:0], dOut);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
