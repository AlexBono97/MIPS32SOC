//  A testbench for testMemDecoder_tb
`timescale 1us/1ns

module testMemDecoder_tb;
    reg [31:0] vAddr;
    reg mWrite;
    reg mRead;
    wire [12:0] pAddr;
    wire [2:0] mEnab;
    wire [1:0] mBank;
    wire iAddr;

  testMemDecoder testMemDecoder0 (
    .vAddr(vAddr),
    .mWrite(mWrite),
    .mRead(mRead),
    .pAddr(pAddr),
    .mEnab(mEnab),
    .mBank(mBank),
    .iAddr(iAddr)
  );

    reg [52:0] patterns[0:55];
    integer i;

    initial begin
      patterns[0] = 53'b00010000000000010000000000000000_0_1_0000000000000_001_00_0;
      patterns[1] = 53'b00010000000000010000000000000001_0_1_0000000000001_001_00_0;
      patterns[2] = 53'b00010000000000010000000000000010_0_1_0000000000010_001_00_0;
      patterns[3] = 53'b00010000000000010000000000000011_0_1_0000000000011_001_00_0;
      patterns[4] = 53'b00010000000000010000000000000000_1_0_0000000000000_001_00_0;
      patterns[5] = 53'b00010000000000010000000000000001_1_0_0000000000001_001_00_0;
      patterns[6] = 53'b00010000000000010000000000000010_1_0_0000000000010_001_00_0;
      patterns[7] = 53'b00010000000000010000000000000011_1_0_0000000000011_001_00_0;
      patterns[8] = 53'b00010000000000001111111111111111_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[9] = 53'b00010000000000001111111111111111_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[10] = 53'b00010000000000010001000000000000_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[11] = 53'b00010000000000010001000000000000_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[12] = 53'b00010000000000010000111111111111_0_1_0111111111111_001_00_0;
      patterns[13] = 53'b00010000000000010000111111111111_1_0_0111111111111_001_00_0;
      patterns[14] = 53'b01111111111111111110111111111100_0_1_1000000000000_001_00_0;
      patterns[15] = 53'b01111111111111111110111111111101_0_1_1000000000001_001_00_0;
      patterns[16] = 53'b01111111111111111110111111111110_0_1_1000000000010_001_00_0;
      patterns[17] = 53'b01111111111111111110111111111111_0_1_1000000000011_001_00_0;
      patterns[18] = 53'b01111111111111111110111111111100_1_0_1000000000000_001_00_0;
      patterns[19] = 53'b01111111111111111110111111111101_1_0_1000000000001_001_00_0;
      patterns[20] = 53'b01111111111111111110111111111110_1_0_1000000000010_001_00_0;
      patterns[21] = 53'b01111111111111111110111111111111_1_0_1000000000011_001_00_0;
      patterns[22] = 53'b01111111111111111110111111111011_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[23] = 53'b01111111111111111110111111111011_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[24] = 53'b01111111111111111111111111111100_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[25] = 53'b01111111111111111111111111111100_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[26] = 53'b01111111111111111111111111111011_0_1_1111111111111_001_00_0;
      patterns[27] = 53'b01111111111111111111111111111011_1_0_1111111111111_001_00_0;
      patterns[28] = 53'b00000000000000001011100000000000_0_1_0000000000000_010_01_0;
      patterns[29] = 53'b00000000000000001011100000000001_0_1_0000000000001_010_01_0;
      patterns[30] = 53'b00000000000000001011100000000010_0_1_0000000000010_010_01_0;
      patterns[31] = 53'b00000000000000001011100000000011_0_1_0000000000011_010_01_0;
      patterns[32] = 53'b00000000000000001011100000000000_1_0_0000000000000_010_01_0;
      patterns[33] = 53'b00000000000000001011100000000001_1_0_0000000000001_010_01_0;
      patterns[34] = 53'b00000000000000001011100000000010_1_0_0000000000010_010_01_0;
      patterns[35] = 53'b00000000000000001011100000000011_1_0_0000000000011_010_01_0;
      patterns[36] = 53'b00000000000000001011011111111111_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[37] = 53'b00000000000000001011011111111111_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[38] = 53'b00000000000000001100101011000000_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[39] = 53'b00000000000000001100101011000000_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[40] = 53'b00000000000000001100101010111111_0_1_1001010111111_010_01_0;
      patterns[41] = 53'b00000000000000001100101010111111_1_0_1001010111111_010_01_0;
      patterns[42] = 53'b11111111111111110000000000000000_0_1_0000000000000_100_10_0;
      patterns[43] = 53'b11111111111111110000000000000001_0_1_0000000000001_100_10_0;
      patterns[44] = 53'b11111111111111110000000000000010_0_1_0000000000010_100_10_0;
      patterns[45] = 53'b11111111111111110000000000000011_0_1_0000000000011_100_10_0;
      patterns[46] = 53'b11111111111111110000000000000000_1_0_0000000000000_100_10_0;
      patterns[47] = 53'b11111111111111110000000000000001_1_0_0000000000001_100_10_0;
      patterns[48] = 53'b11111111111111110000000000000010_1_0_0000000000010_100_10_0;
      patterns[49] = 53'b11111111111111110000000000000011_1_0_0000000000011_100_10_0;
      patterns[50] = 53'b11111111111111101111111111111111_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[51] = 53'b11111111111111101111111111111111_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[52] = 53'b11111111111111110000000000010000_1_0_xxxxxxxxxxxxx_000_xx_1;
      patterns[53] = 53'b11111111111111110000000000010000_0_1_xxxxxxxxxxxxx_000_xx_1;
      patterns[54] = 53'b11111111111111110000000000001111_0_1_0000000001111_100_10_0;
      patterns[55] = 53'b11111111111111110000000000001111_1_0_0000000001111_100_10_0;

      for (i = 0; i < 56; i = i + 1)
      begin
        vAddr = patterns[i][52:21];
        mWrite = patterns[i][20];
        mRead = patterns[i][19];
        #10;
        if (patterns[i][18:6] !== 13'hx)
        begin
          if (pAddr !== patterns[i][18:6])
          begin
            $display("%d:pAddr: (assertion error). Expected %h, found %h", i, patterns[i][18:6], pAddr);
            $finish;
          end
        end
        if (patterns[i][5:3] !== 3'hx)
        begin
          if (mEnab !== patterns[i][5:3])
          begin
            $display("%d:mEnab: (assertion error). Expected %h, found %h", i, patterns[i][5:3], mEnab);
            $finish;
          end
        end
        if (patterns[i][2:1] !== 2'hx)
        begin
          if (mBank !== patterns[i][2:1])
          begin
            $display("%d:mBank: (assertion error). Expected %h, found %h", i, patterns[i][2:1], mBank);
            $finish;
          end
        end
        if (patterns[i][0] !== 1'hx)
        begin
          if (iAddr !== patterns[i][0])
          begin
            $display("%d:iAddr: (assertion error). Expected %h, found %h", i, patterns[i][0], iAddr);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
